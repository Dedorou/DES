module encrypt_tb();

reg clk = 0;
reg [0 : 63] data_in;
wire [0 : 63] data_out;
reg [0 : 47] key;
reg mux, load;
wire ready;

parameter clk_period = 100;

always #(clk_period/2) clk=~clk;

encryption_block encr (clk, 1'b0, data_in, key, 1'b0, mux, load, data_out);	

initial begin 

mux = 0;
load = 0;
data_in = 64'b0000000011100000000011101110000000001110111011101110111000000000;
#clk_period;
#clk_period;
#clk_period;
load <= 1;
#clk_period;
mux <= 1;
key <= 64'b000100000000000011101100001100000010100011000011;
#clk_period;
key <= 64'b010100001010110011010000011100100010000101000101;

#clk_period;
key <= 64'b010101001110110000000010101000101000000110001010;
#clk_period;
key <= 64'b011000101010010100000110010001000011011100000011;
#clk_period;
key <= 64'b011010001000010000000111011111100000000001101000;
#clk_period;
key <= 64'b011000011000000000111010010000001101100101001010;
#clk_period;
key <= 64'b101001001000000010110010000001001011010000111000;
#clk_period;
key <= 64'b101101100000101000010010111010010001110001100000;
#clk_period;
key <= 64'b001000000101101101000011010010111101001000100000;
#clk_period;
key <= 64'b001000010111000101000101100100000100110100101000;
#clk_period;
key <= 64'b000000010100010111010001100010000001101000010100;
#clk_period;
key <= 64'b010101010100000110110001110100010110001010110000;
#clk_period;
key <= 64'b100101111000000110000001001100010000101000001001;
#clk_period;
key <= 64'b000110110000001010000111100100100011000000010110;
#clk_period;
key <= 64'b001110010001000010001100001001010010001110100100;
#clk_period;
key <= 64'b010000010011110010001000000001100110001010000001;
#clk_period;
#clk_period;

end

endmodule 




/*
64'b000100000000000011101100001100000010100011000011


64'b010100001010110011010000011100100010000101000101

64'b010101001110110000000010101000101000000110001010

64'b011000101010010100000110010001000011011100000011

64'b011010001000010000000111011111100000000001101000

64'b011000011000000000111010010000001101100101001010

64'b101001001000000010110010000001001011010000111000

64'b101101100000101000010010111010010001110001100000

64'b001000000101101101000011010010111101001000100000

64'b001000010111000101000101100100000100110100101000

64'b000000010100010111010001100010000001101000010100

64'b010101010100000110110001110100010110001010110000

64'b100101111000000110000001001100010000101000001001

64'b000110110000001010000111100100100011000000010110

64'b001110010001000010001100001001010010001110100100

64'b010000010011110010001000000001100110001010000001
*/










