module crypt_block
(input [0 : 63] data_in)

endmodule